/*
 * Copyright 2019 ISP RAS (http://www.ispras.ru)
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     http://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 */

// IEEE Std 1800-2012
//   16. Assertions
//    16.9 Sequence operations
//     16.9.5 AND operation

// ! TYPE: POSITIVE

module test;

reg te1, te2, te3, te4, te5;

sequence seq1;
  (te1 ##2 te2) and (te3 ##2 te4 ##2 te5);
endsequence

sequence seq2;
  (te1 ##[1:5] te2) and (te3 ##2 te4 ##2 te5);
endsequence

endmodule
