/*
 * Copyright 2018 ISP RAS (http://www.ispras.ru)
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     http://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 */

// IEEE Std 1364-2005
//   6. Expressions
//     6.1 Continuous assignments
//       6.1.2 The continuous assignment statement
//         The following is an example of a continuous assignment to a net that
//         has been previously declared

module test;
  reg enable;
  wire  mynet;
  assign (strong1, pull0) mynet = enable;
endmodule
