/*
 * Copyright 2018 ISP RAS (http://www.ispras.ru)
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     http://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 */

// IEEE Std 1364-2005
//   5. Expressions
//    5.1 Operators
//      5.1.7 Relational operators
//        Table 5-10 - Definitions of relational operators

module test;

  integer a, b, c;

  initial begin
    c = a < b;  // a less than b
    c = a > b;  // a greater than b
    c = a <= b; // a less than or equal to b
    c = a >= b; // a greater than or equal to b
  end
endmodule
