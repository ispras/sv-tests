/*
 * Copyright 2018-2024 ISP RAS (http://www.ispras.ru)
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     http://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 */

// IEEE Std 1364-2005
//   15. Timing checks
//     15.2 Timing checks using a stability window
//       15.2.3 $setuphold
//         The $setuphold timing check combines the functionality of the $setup and $hold timing
//         checks into a single timing check.

module test(clk, data);
  input clk, data;

  specify
    specparam tSU = 1.5, tHLD = 2.1;
    $setuphold (posedge clk, data, tSU, tHLD);
    // is equivalent in functionality to the following, if tSU and tHLD are not negative
    $setup (data, posedge clk, tSU);
    $hold (posedge clk, data, tHLD);
  endspecify
endmodule
