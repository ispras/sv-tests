/*
 * Copyright 2018 ISP RAS (http://www.ispras.ru)
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     http://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 */

// IEEE Std 1364-2005
//   4. Data types
//    4.9 Arrays
//      4.9.3 Memories
//        4.9.3.1 Array examples
//          4.9.3.1.1 Array declarations
module test;
  reg [7:0] mema[0:255];   // declares a memory mema of 256 8-bit
                           // registers. The indices are 0 to 255
  reg arrayb[7:0][0:255];  // declare a two-dimensional array of
                           // one bit registers
  wire w_array[7:0][5:0];  // declare array of wires
  integer inta[1:64];      // an array of 64 integer values
  time chng_hist[1:1000];  // an array of 1000 time values
  integer t_index;
endmodule
