/*
 * Copyright 2018 ISP RAS (http://www.ispras.ru)
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     http://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 */

// IEEE Std 1364-2005
//   12. Hierarchical structures
//     12.3 Ports
//       12.3.6 Connecting module instance ports by name
//         Multiple module instance port connections are not allowed, e.g., the following example is
//         illegal. This example shows illegal port connections.

// ! TYPE: VARYING

module test;

`ifdef NEGATIVE_TEST
  a ia (.i (a), .i (b),  // illegal connection of input port twice.
        .o (c), .o (d),  // illegal connection of output port twice.
        .e (e), .e (f)); // illegal connection of inout port twice.
`endif
endmodule
